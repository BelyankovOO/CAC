module instructionmemory(input [31:0] addr, output reg [31:0] com);

always @(addr)
	case(addr)
		32'h00000000: com <= 32'b001000_00000_10000_0000000000000111; //addi r16 r0 7
		32'h00000004: com <= 32'b101011_00000_10000_0000000000000001; //sw M[1+r0] <- r16

		32'h00000008: com <= 32'b100011_00000_10011_0000000000000001; //lw M[1+r0] -> r19
		32'h0000000c: com <= 32'b000000_10011_00100_00011_00000_100000; //add r3 = r19 + r4 

		//32'h00000000: com <= 32'b001000_00000_10011_0000000000000100; //addi r19 = r0 + 4
		//32'h00000004: com <= 32'b000000_10011_10001_00001_00000_100000; //add r1 = r19 + r17
		//32'h00000008: com <= 32'b000000_00001_10011_00010_00000_100000; //add r2 = r1 + r19
        
		//32'h00000000: com = 32'b001000_00000_10001_0000000000000011; //addi r17 = r0 + 3
		//32'h00000004: com = 32'b001000_10001_10010_0000000000000001; //addi r18 = r17 + 1
		//32'h00000008: com = 32'b001000_10001_10011_0000000000000010; //addi r19 = r17 + 2

		//32'h00000008: com = 32'b000100_10000_10001_0000000000001100; //beq //24
		//32'h0000000c: com = 32'b001000_10000_10000_0000000000000001; //addi
		//32'h00000010: com = 32'b000100_10000_10001_0000000000001000; //beq //16
		//32'h00000014: com = 32'b001000_10000_10000_0000000000000001; //addi
		//32'h00000018: com = 32'b000100_10000_10001_0000000000000100; //beq //8
		//32'h0000001c: com = 32'b001000_10000_10000_0000000000000001; //addi

		//32'h00000020: com = 32'b001000_00000_10011_0000000000001111; //addi
		//32'h00000024: com = 32'b000010_00000000000000000000000100;//j 4

		//32'h00000004: com <= 32'b001000_00000_10000_0000000000000011; //addi s0 0 c

		default: com <= 32'b111111_00000_00000_0000000000000000; //noop
	endcase 
	
endmodule		
