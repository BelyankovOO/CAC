module instructionmemory(input [31:0] addr, output reg [31:0] com);

always @(addr)
	case(addr)
		//32'h00000000: com <= 32'b001000_00000_10000_0000000000000111; //addi s0 0 c
		//32'h00000004: com <= 32'b101011_00000_10000_0000000000000001; //sw s0 1
		//32'h00000008: com <= 32'b100011_00000_10010_0000000000000001; //lw s2 1
		//32'h0000000c: com <= 32'b100011_00000_10001_0000000000000001; //lw s1 1
		//32'h00000010: com <= 32'b000000_10010_10001_10011_00000_100000; //add s2 s1 s0
        
		32'h00000000: com <= 32'b001000_00000_10001_0000000000000011; //addi s1 0 c

		32'h00000004: com <= 32'b001000_10000_10000_0000000000000001; //addi s0 s0 c
		32'h00000008: com <= 32'b000100_10000_10001_0000000000100000; //beq
		32'h0000000c: com <= 32'b001000_10000_10000_0000000000000001; //addi
		32'h00000010: com <= 32'b000100_10000_10001_0000000000100000; //beq
		32'h00000014: com <= 32'b001000_10000_10000_0000000000000001; //addi
		32'h00000018: com <= 32'b000100_10000_10001_0000000000100000; //beq
		32'h0000001c: com <= 32'b001000_10000_10000_0000000000000001; //addi

		32'h00000020: com <= 32'b001000_00000_10011_0000000000001111; //addi

		//32'h00000004: com <= 32'b001000_00000_10000_0000000000000011; //addi s0 0 c

		default: com <= 0;
	endcase 
	
endmodule		
